Project1	project	Next Generation Analysis Tools	bioinfo	Bioinformatics Team
skhuri	user	Sawsan Khuri	bioinfo	Bioinformatics Team
Project2	project	Next Generation Data Analysis	nextgen	Next Generation Sequencing
yedwards	user	Yvonne Edwards	nextgen	Next Generation Sequencing
dhedges	user	Dale Hedges	nextgen	Next Generation Sequencing

